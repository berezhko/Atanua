module not6 (
    input [5:0] a,
    output reg [5:0] out
);

assign out = ~a;

endmodule
