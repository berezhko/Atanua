module myor (
    input wire a,
    input wire b,
    output reg out
);

assign out = a | b;

endmodule
